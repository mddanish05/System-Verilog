interface intf;
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic carry;
endinterface
